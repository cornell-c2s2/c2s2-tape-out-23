module logo_svg ();
endmodule