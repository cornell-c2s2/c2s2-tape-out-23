// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_project_wrapper
 *
 * This wrapper enumerates all of the pins available to the
 * user for the user project.
 *
 * An example user project is provided in this wrapper.  The
 * example should be removed and replaced with the actual
 * user project.
 *
 *-------------------------------------------------------------
 */

module user_project_wrapper #(
    parameter BITS = 32
) (
`ifdef USE_POWER_PINS
    inout vdda1,	// User area 1 3.3V supply
    inout vdda2,	// User area 2 3.3V supply
    inout vssa1,	// User area 1 analog ground
    inout vssa2,	// User area 2 analog ground
    inout vccd1,	// User area 1 1.8V supply
    inout vccd2,	// User area 2 1.8v supply
    inout vssd1,	// User area 1 digital ground
    inout vssd2,	// User area 2 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // Analog (direct connection to GPIO pad---use with caution)
    // Note that analog I/O is not available on the 7 lowest-numbered
    // GPIO pads, and so the analog_io indexing is offset from the
    // GPIO indexing by 7 (also upper 2 GPIOs do not have analog_io).
    inout [`MPRJ_IO_PADS-10:0] analog_io,

    // Independent clock (on independent integer divider)
    input   user_clock2,

    // User maskable interrupt signals
    output [2:0] user_irq
);

/*--------------------------------------*/
/* User project is instantiated  here   */
/*--------------------------------------*/

FFTSPIInterconnectRTL fft_spi
(
`ifdef USE_POWER_PINS
    .vccd1(vccd1),	// User area 1 1.8V supply
    .vssd1(vssd1),	// User area 1 digital ground
`endif
  .clk            ( wb_clk_i    ),
  .reset          ( wb_rst_i    ),

  // Inputs

  .minion_sclk    ( io_in[11]   ),
  .minion_sclk_2  ( io_in[15]   ),
  .minion_sclk_3  ( io_in[19]   ),
  .minion_mosi    ( io_in[10]   ),
  .minion_mosi_2  ( io_in[14]   ),
  .minion_mosi_3  ( io_in[18]   ),
  .minion_cs      ( io_in[9]    ),
  .minion_cs_2    ( io_in[13]   ),
  .minion_cs_3    ( io_in[17]   ),

  .master_miso    ( io_in[22]   ),

  // Outputs

  .adapter_parity ( io_out[7]   ),
  .minion_parity  ( io_out[8]   ),
  .minion_miso    ( io_out[12]  ),
  .minion_miso_2  ( io_out[16]  ),
  .minion_miso_3  ( io_out[20]  ),
  .master_cs      ( io_out[21]  ),
  .master_mosi    ( io_out[23]  ),
  .master_sclk    ( io_out[24]  ),

  // Output Enables


  .io_oeb         (  )
);

assign io_oeb[24:7] = 18'b001001110111011100; // Will Fed up the io_oeb due to sleep deprivation so assigning it here so we 
//don't need to wait like 16 hours to push through the flow again. 
endmodule	// user_project_wrapper

`default_nettype wire